`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Dependencies: 
//
// Revision 3.0

// Additional Comments: for Z80 bus
//
//////////////////////////////////////////////////////////////////////////////////
module main(
				//CPU
				a_cpu,
				d_cpu,
				wr_cpu,rd_cpu,io_req_cpu,reset_cpu,clk_cpu,
				iei,ieo,
				m1_cpu,
				int_cpu,
				nmi_cpu,
				mem_req_cpu,
				rfsh_cpu,
				halt_cpu,
				wait_cpu,
				bus_req_cpu,
				bus_ack_cpu,
				reserved_cpu,
				
				watchdog,
				
				//OSC
				clk_scan, 
				
				//RAM
				a_ram,
				d_ram,
				oe_ram,
				wr_ram,
				cs_ram_out,
				cs_ram_in,
				
			
				//TAP 1
				tdo_1,
				tck_1,
				tms_1,
				trst_1,
				tdi_1,
				fail_1,

				//TAP 2
				tdo_2,
				tck_2,
				tms_2,
				trst_2,
				tdi_2,
				fail_2,

				//GPIO
				gpio,
				
				//DEBUG
				debug,
				
				// start/stop/sts front panel
				start,
						// synthesis attribute PULLUP of start is“TRUE”;
				stop,
						// synthesis attribute PULLUP of stop is“TRUE”;
				pass,
				fail,
	
				// UUT pwr control
				uut_pwr_on_1,
				uut_pwr_on_2,
				uut_pwr_fail_1,	
				uut_pwr_fail_2,		
	
				//pwr_good
				//pwr_good,
	
				//I2C
				sda,
				scl,
				
				rsv_16
								
				);
	
	// CPU
	input [15:0] a_cpu;
	inout [7:0] d_cpu; 
   input wr_cpu;
	input reset_cpu;
	input rd_cpu;
   input io_req_cpu;
	input clk_cpu;
	input iei;
	input	ieo;
	input m1_cpu;
	output int_cpu;
	assign int_cpu = 1'bz;  //temporarily
	output nmi_cpu;
	assign nmi_cpu = 1'bz;  //temporarily
	input mem_req_cpu;
	input rfsh_cpu;
	input	halt_cpu;
	output wait_cpu;
	assign wait_cpu = 1'bz; //temporarily
	input bus_req_cpu;	//CS: not sure , check !
	input bus_ack_cpu;	//CS: not sure , check !
	input [7:0] reserved_cpu;

	input watchdog;
		// synthesis attribute PULLUP of watchdog is TRUE;
		
	//RAM
   output oe_ram;
   output wr_ram;
	output cs_ram_out;
	output cs_ram_in;
	assign cs_ram_in = 1'b1; //temporarily

   output [23:0] a_ram;
		// synthesis attribute PULLUP of a_ram is“TRUE”;
   inout [7:0] d_ram;
		// synthesis attribute PULLUP of d_ram is“TRUE”;


	// GPIO
	inout [3:0] gpio;
	
	// tap 1
   output tdo_1;
	output tms_1;
   output tck_1;
   output trst_1;
	input tdi_1;
	output fail_1;
	//assign fail_1 = 1'bz;  //temporarily

	// tap 2
   output tdo_2;
	output tms_2;
   output tck_2;
   output trst_2;
	input tdi_2;
	output fail_2;
	assign fail_2 = 1'bz;  //temporarily	
	
	// OSC
   input clk_scan;
	 
	
	//rsv
	input rsv_16;	 // 1 hz clock
	 
	 
	// debug
	output [7:0] debug;
	//assign debug[7:3] = 6'h00;  //temporarily
	//assign debug[2] = !tck_1; //blue
	//assign debug[0] = !fail_1; //rsv_16; //red

	// start/stop/sts front panel
	input start;
	input stop;
	output pass;
	output fail;	

	
	// UUT pwr control
	// use fail_any_chain for PWR off !
	output uut_pwr_on_1;
	assign uut_pwr_on_1 = 1'bz; //temporarily
	
	output uut_pwr_on_2;
	assign uut_pwr_on_2 = 1'bz; //temporarily
	
	output uut_pwr_fail_1;	
	assign uut_pwr_fail_1 = 1'bz; //temporarily
	output uut_pwr_fail_2;		
	assign uut_pwr_fail_2 = 1'bz; //temporarily
	
	// watchdog
	//input watchdog;
	
	//pwr_good
	//input pwr_good;
	
	//I2C
	inout sda;
	// synthesis attribute FLOAT of sda is“TRUE”;
	inout scl;
	// synthesis attribute FLOAT of scl is“TRUE”;

/////////////////////////////////////////////////////////////////////////////////////////

	`include "parameters.v"
	

	wire data_write_strobe;
	wire [63:0] gpo_rf;
	wire [215:0] gpi_rf;
	
	reg_file_z80 rf (
		.a_cpu(a_cpu[7:0]), 
		.d_cpu(d_cpu), 
		.wr_cpu(wr_cpu), 
		.rd_cpu(rd_cpu),
		.io_req_cpu(io_req_cpu), 
		.reset_cpu(reset_cpu),
		.clk_cpu(clk_cpu),
		.general_purpose_out(gpo_rf[63:0]),		//  [7:0] 80h -> data channel write access
														//	[31:8] 83-81h -> ram address
														// [39:32] 84h -> command channel
														// [47:40] 8Bh -> signal path
														// [55:48] 8Ch -> frequency
														// [63:56] 89 -> test start/stop (55/AA)
														
		.general_purpose_in(gpi_rf[215:0]),		//  [7:0] 80h -> data channel read access
														// [31:8] 87-85h -> for debug: RAM address generated by executor
														
														// [34:32] 88h -> for debug: selected bit address generated by executor
														// [35] 88h -> for debug: bit data of selected bit
														
														// [39:32] 88h -> fail_1,exp_1,tdi_1,mask_1
														
														// [47:40] 89h -> executor state
														// [55:48] 8Ah -> tap states
														// [87:56] 8F-8Ch -> bits processed chain 1
														// [119:88]	93-90 -> sxr_length_chain_1
														// [135:120] 95-94 -> step id
														// [143:136] 96 -> vec_state_1
														// [175:144] 9A-97 -> bits processed chain 2
														// [207:176] 9E-9B -> sxr_length_chain_2
														// [215:208] 9F -> vec_state_2
		.data_write_strobe(data_write_strobe) // L on write access to 80h (data channel)
	);

	
	
	
	
	wire [7:0] path;
	assign path = gpo_rf[47:40];
	
	wire [7:0] command;
	assign command = gpo_rf[39:32]; // write to 84h


	// RAM signals routing
	wire [23:0] a_ram_rf;
	assign a_ram_rf = gpo_rf[31:8]; //rf write address 83-81h 
	wire [23:0] a_ram_ex;
	reg [23:0] a_ram;
	assign gpi_rf[31:8] = a_ram; // rf may read any time at 87-85h from a_ram
	
	wire [7:0] d_ram_rf;
	assign d_ram_rf = gpo_rf[7:0];
	wire [7:0] d_ram_ex;
	assign d_ram_ex = d_ram;	// ex always reads data from RAM
	assign gpi_rf[7:0] = d_ram; // rf may read any time at 80h from d_ram;
	
	// address
	// source is rf or ex
	always @*
		begin
			case (path[3:2])
				2'b00	: a_ram = a_ram_rf; // rf drives adr in RAM // write adr 83-81h
				2'b01 : a_ram = a_ram_ex; // ex reads from RAM
				default : a_ram = 8'hzz; // on reset or pwr-up //  pull-ups internally
			endcase
		end
		

	// data
	// source is rf or output RAM
	reg wr_ram;
	reg oe_ram;
	reg cs_ram_out;
	always @*
		begin
			case (path[1:0])
				2'b00 : 	// rf writes in RAM
					begin
						wr_ram = data_write_strobe; // on write to rf 80h
						oe_ram = 1'b1; // RAM read forbidden
						cs_ram_out = 1'b0; // CS: should depend on ram address
					end

				2'b01 : 	// reading from RAM
					begin
						wr_ram = 1'b1; // RAM write forbidden
						oe_ram = 1'b0;
						cs_ram_out = 1'b0; // CS: should depend on ram address
					end
				
				default : // on reset or pwr-up 
					begin 
						wr_ram = 1'b1; 
						oe_ram = 1'b1; 
						cs_ram_out = 1'b1; 						
					end
			endcase
		end
		
		assign d_ram = oe_ram ? d_ram_rf : 8'hzz; // drive data to RAM if oe_ram=1 , else release d_ram
		

	clk_divider cd (
		.clk_in(clk_scan),
		.clk_out(clk_test),
		.reset(reset_cpu),
		.scale(gpo_rf[55:48]) //8C
    );


	// STS LED and debug
	reg step_mode;
	wire clk_led;
	wire clk_debouncer;
	always @*
		begin
			case (command[3:0])
				tck_step	:	step_mode <= clk_led;
				sxr_step	:	step_mode <= clk_debouncer; // fast led flashing derived from debouncer clock
				default	:	step_mode <= 1;
			endcase
		end
		
	reg [7:0] debug;
	wire test_running;
	wire led;
	wire tap_ready;
	always @*
		begin
			casex ({path[3:0],test_running})
				5'b0001x	: 	begin
									debug[1] = rsv_16; // yellow LED flashes to indicate RAM read/debug mode
									debug[2] = 1'b1;   // blue LED off
								end
				5'b01011	: 	begin
									debug[1] = 1'b1;   // yellow LED off
									debug[2] = rsv_16; // blue LED flashes to indicate executor mode idle
								end
				5'b01010	: 	begin
									debug[1] = step_mode; // yellow flashes fast on sxr_step_width, slow on tck_step_width
									debug[2] = 1'b0; // blue LED on to indicate executor is running
									debug[0] = !fail; // red flashes on fail
									debug[3] = clk_test;
									//debug[4] = clk_test;
								end
				5'b0000x	: 	begin
									debug[1] = 1'b0;   // yellow LED on to indicate RAM write mode
									debug[2] = 1'b1;   // blue LED off
								end
				default	: debug = 8'hFF;   // all LED off after reset or pwr up //
			endcase
		end
		
		
	prescaler ps (
		.clk(clk_cpu),
		.qf(clk_debouncer),	// fast flashing leds	// updated on posedge of cpu_clk
		.qg(clk_led)			// slow flashing leds  	// updated on posedge of cpu_clk
	);
	
	
	wire [7:0] strt_stop;
	assign strt_stop = gpo_rf[63:56]; //98  // updated on posedge of cpu_clk
	reg start_rf;
	reg stop_rf;
	always @(negedge clk_cpu)
		begin
			case (strt_stop)
				8'hAA		: 	begin	// stop test
									start_rf <= 1;
									stop_rf <= 0;
								end
				8'h55		: 	begin	// start test
									start_rf <= 0;
									stop_rf <= 1;
								end
				default	: 	begin
									start_rf <= 1;
									stop_rf <= 1;
								end
			endcase
		end
				
	debouncer db_start (
		.out(start_db),  // L-active  // updated on nededge of clk
		.in(start),  // L-active  from start button front panel
		.clk(clk_debouncer)  
	);

	assign start_x = (start_rf & start_db); 	// collect start signals here  //start_x updated on negedge clk_cpu
	
	


	debouncer db_stop (
		.out(stop_db),  // L-active  // updated on nededge of clk
		.in(stop),  // L-active  from stop button front panel
		.clk(clk_debouncer)
	);

	assign stop_x = (stop_rf & stop_db);	// collect stop signals here  //stop_x updated on negedge clk_cpu


	
	
	wire [31:0] bits_processed_chain_1;
	wire [31:0] bits_processed_chain_2;	
	wire [31:0] sxr_length_chain_1;
	wire [31:0] sxr_length_chain_2;	
	wire [15:0] step_id;
	
	wire [7:0] vec_state_1;	
	wire [7:0] vec_state_2;
	
	executor ex (
		.reset(reset_cpu),
		.start(start_x),	// L-active
		.stop(stop_x),	// L-active
		//.active(test_running),	//ouput; address controlled by executor ex // L active
		.start_addr(a_ram_rf), 			//driven by register file //83-81h
		.ram_addr(a_ram_ex), 			//drives output RAM address (if executor control selected)
		.ram_data(d_ram_ex),				//driven by d_ram
		//.selected_bit(gpi_rf[34:32]),	//outputs address of selected bit of RAM data
		//.bit_data(gpi_rf[36]),			//outputs selected bit data
		.tdi_1(tdi_1),
		.tdi_2(tdi_2),
		.tdo_1(tdo_1),
		.tdo_2(tdo_2),
		.tms_1(tms_1),
		.tms_2(tms_2),
		.tck_1(tck_1),
		.tck_2(tck_2),
		.trst_1(trst_1),
		.trst_2(trst_2),
		.fail_1(fail_1),  // H - active
		.fail_2(fail_2),
		.fail_any_chain(fail_any_chain), // H-active (when ex in test_fail)
		.step_id(step_id),
		.pass(pass),
		.mask_1(mask_1),
		.mask_2(mask_2),
		.exp_1(exp_1),
		.exp_2(exp_2),		
		//.clk_cpu(clk_cpu),
		.clk(clk_test), // (rsv_16),		//CS: drive clk_tap via on board osc and prescaler
		//.mode(gpo_rf[39:32]),	//rf command channel output // 84h
		.mode(command),		//halt executor on FFh , start on 10h
		.exec_state(gpi_rf[47:40]),  //read from 89h
		.run(test_running),  // run is L-active
		.debug(gpi_rf[55:48]),  // read from 8A
		//.led(led),
		.bits_processed_chain_1(bits_processed_chain_1),
		.bits_processed_chain_2(bits_processed_chain_2),
		.sxr_length_chain_1(sxr_length_chain_1),
		.sxr_length_chain_2(sxr_length_chain_2),
		//.bit_no_1(bit_no_1),
		//.bit_no_2(bit_no_2),
		.tap_ready(tap_ready),
		.vec_state_1(vec_state_1),
		.vec_state_2(vec_state_2)
	);

	// [143:136] 96 -> vec_state_1 (from tc)
	// [151:144] 97 -> bit [7:5]=0, [4:0] bit_no_2 from tc
	assign gpi_rf[143:136] = vec_state_1; // 96
	assign gpi_rf[215:208] = vec_state_2; // 9F



	assign fail = fail_any_chain & clk_debouncer;

	//	wire [31:0] bits_processed_chain_1_dec;
	//	assign bits_processed_chain_1_dec[31:0] = bits_processed_chain_1[31:0] -1; //on fail bits_processed_chain_1 is one bit ahead, so subtract 1

		assign gpi_rf[63:56] = bits_processed_chain_1[7:0];  // 8C
		assign gpi_rf[71:64] = bits_processed_chain_1[15:8];
		assign gpi_rf[79:72] = bits_processed_chain_1[23:16];
		assign gpi_rf[87:80] = bits_processed_chain_1[31:24];	// 8F	

		assign gpi_rf[95:88]   = sxr_length_chain_1[7:0];  	// 90
		assign gpi_rf[103:96]  = sxr_length_chain_1[15:8];
		assign gpi_rf[111:104] = sxr_length_chain_1[23:16];
		assign gpi_rf[119:112] = sxr_length_chain_1[31:24];	// 93
		
		assign gpi_rf[135:120] = step_id[15:0];	// 95-94
		
		assign gpi_rf[175:144] = bits_processed_chain_2[31:0]; // 9A-97
		assign gpi_rf[207:176] = sxr_length_chain_2[31:0]; 	// 9E-9B

		assign gpi_rf[39:32]	= {fail_2,exp_2,tdi_2,mask_2,fail_1,exp_1,tdi_1,mask_1}; //88

endmodule


//////O L D///////////////////////////////////////////////////////////////////////////////////////////////
/*
	wire [23:0] a_ram_executor;
	wire run;
	reg [7:0] mode_ex;
	//assign addr_by_rf_or_ex = 1'b1;
	executor ex (
		.active(addr_by_rf_or_ex),	//ouput; address controlled by executor ex // L active
		.start_addr(gpo_rf[31:8]), 	//driven by register file //83-81h
		.ram_addr(a_ram_executor), //drives output RAM address (if executor control selected)
		.ram_data(d_ram),		//driven by output RAM
		.selected_bit(gpi_rf[34:32]),	//outputs address of selected bit of RAM data
		.bit_data(gpi_rf[36]),			//outputs selected bit data
		.tdo_1(tdo_1),
		.tdo_2(tdo_2),
		.tms_1(tms_1),
		.tms_2(tms_2),
		.tck_1(tck_1),
		.tck_2(tck_2),
		.trst_1(trst_1),
		.trst_2(trst_2),
		.fail_1(fail_1),
		.fail_2(fail_2),
		.clk_cpu(clk_cpu),
		.clk_tap(rsv_16),		//CS: drive clk_tap via on board osc and prescaler
		//.mode(gpo_rf[39:32]),	//rf command channel output // 84h
		.mode(mode_ex),	//made by mode decoder
		.exec_state(gpi_rf[47:40]),  //89h
		.run(run),
		.debug(gpi_rf[55:48])
	);
	
	assign gpi_rf[31:8] = a_ram_executor;	//for debugging executor 87-85h
	assign gpi_rf[39:37] = 3'b000;
	assign gpi_rf[35] = 1'b0;

	// output RAM signal mapping begin
	assign a_ram = addr_by_rf_or_ex ? gpo_rf[31:8] : a_ram_executor; // gpo[31:8] -> 83-81h
	assign gpi_rf[7:0] = d_ram;   //read from 80h
	
	//assign d_ram = data_write_strobe ? 8'hzz : gpo_rf[7:0];  //write to 80h	
	reg [7:0] d_ram_rf;
	reg wr_ram;
	always @*
		begin
			case (gpo_rf[39:32])  //mode (written in cmd channel 84h)
				8'hFF	:	begin
								d_ram_rf = gpo_rf[7:0];  //write to 80h
								wr_ram = data_write_strobe;
								mode_ex = 8'hFF;	// makes ex idling
							end

				8'h80	:	begin
								d_ram_rf = 8'hzz;
								wr_ram = 1'b1;
								mode_ex = 8'h80;	// gives ex a GO
							end

				default : 
							begin
								d_ram_rf = 8'hzz;
								wr_ram = 1'b1;
								mode_ex = 8'hFF;	// makes ex idling								
							end
			endcase
		end
				
	//assign d_ram = data_write_strobe ? 8'hzz : gpo_rf[7:0];  //write to 80h	
	assign d_ram = d_ram_rf;  //write to 80h	

	assign oe_ram = (addr_by_rf_or_ex & data_read_strobe);
	//assign wr_ram = data_write_strobe; //CS: combine with addr_by_rf_or_ex ?

	reg cs_ram_out;
	always @*	// make CS signal
		begin
			if (a_ram <= ram_top) cs_ram_out <= 1'b0;
			else cs_ram_out <= 1'b1;
		end
	// output RAM signal mapping end		
		

	assign gpio[3:0] = 4'b0000; // temporarily
	//assign gpio[1] = addr_by_rf_or_ex;
	assign debug[1] = addr_by_rf_or_ex ? rsv_16 : 1'b0; // yellow LED flashes in debug mode / on when exector active
endmodule
*/