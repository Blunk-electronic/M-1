`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Dependencies: 
//
// Revision 3.0

// Additional Comments: for Z80 bus
//
//////////////////////////////////////////////////////////////////////////////////
module tdo_gen(a_cpu,d_cpu,wr_cpu,rd_cpu,io_req_cpu,reset_cpu,clk_cpu,
				clk_scan, // driven by tdi_reader
				oe_ram_drv,a_ram,d_ram_drv,wr_ram_drv_exp_mask,cs_ram,
				tdo_gen,
				tck_gen,
				tms_gen,
				trst_gen,state,tdo_en,
				gpio_a,
				gpio_b,
				gpio_c,
				dmux_sel
				);
	
	// cpu begin			
	input [15:0] a_cpu;
	//	 inout [7:0] reserved;
	inout [7:0] d_cpu;
    input wr_cpu;
	input reset_cpu;
	input rd_cpu;
    input io_req_cpu;
	input clk_cpu;
	// cpu end

	// ram out
    output oe_ram_drv;
	output cs_ram;
    output [23:3] a_ram;
    inout [7:0] d_ram_drv;
    output wr_ram_drv_exp_mask;
	 
	// ram in ?

	// gpio
	input [7:0] gpio_a;
	//input [7:3] gpio_b;	// tdi,dio//	input [0:0] gpio_b;	// tdi,dio
	output [7:0] gpio_b; // yel,blue led
	input [7:0] gpio_c;	// pwr, dac
	
	// tap 
   output tdo_gen;
	output tdo_en;
   output tck_gen;
   output tms_gen;
	output trst_gen;

	// clk local
   input clk_scan;  // driven by tdi_reader
	 
	// debug
	output [3:0] state;
	output [2:0] dmux_sel;
	

	// internal begin
//	wire [23:0] a_ag;
//	wire [23:0] adr_rf;
//	wire [23:0] start_adr_rf;
//	wire [23:0] len_rf;	
//	wire [7:0] dat_rf;	
//	wire [7:0] d_mux;
//	wire [7:0] low_level_ctrl;
//	wire [23:0] mode_rf;

//	reg tms_gen;
//	reg tck_gen;
//	reg tdo_en;
//	reg tdo_2state;

//	wire tms_tsg;
//	wire tck_tsg;
//	wire tdo_dmux;
//	wire tdo_req;

	parameter ram_top = 19'hFFFFF;	// top address of output RAM HM628512 (7FFFFh)

	wire data_write_strobe;
	wire data_read_strobe;	
	wire [39:0] gpo;
	wire [55:0] gpi;

	reg_file_z80 rf (
		.a_cpu(a_cpu), 
		.d_cpu(d_cpu), 
		.wr_cpu(wr_cpu), 
		.rd_cpu(rd_cpu),
		.io_req_cpu(io_req_cpu), 
		.reset_cpu(reset_cpu),
		.clk_cpu(clk_cpu),
		.general_purpose_out(gpo[39:0]),		//  [7:0] 80h -> data channel write access
														//	[31:8] 83-81h -> output ram address channel
														// [39:32] 84h -> command channel
														
		.general_purpose_in(gpi[55:0]),		//  [7:0] 80h -> data channel read access
														// [31:8] 87-85h -> for debug: RAM address generated by executor
														// [34:32] 88h -> for debug: selected bit address generated by executor
														// [35] 88h -> for debug: bit data of selected bit
														// [47:40] 89h -> executor state
		.data_write_strobe(data_write_strobe), // L on write access to 80h (data channel)
		.data_read_strobe(data_read_strobe)  	// L on read access to 80h (data channel)
	);


	//wire [15:0] command;
	//command_decoder cd (
	//	.data_in(gpo[39:32]),		// 84h
	//	.cmd_out(command[15:0])		// H active , after reset all command lines drive L  // updated on posedge of cpu_clk
	//);

	//assign addr_by_rf_or_ex = 1'b1;	// address controlled by executor ex // L active
	wire [23:0] a_ram_executor;
	wire run;
	//assign addr_by_rf_or_ex = 1'b1;
	executor ex (
		.active(addr_by_rf_or_ex),	//ouput; address controlled by executor ex // L active
		.start_addr(gpo[31:8]), 	//driven by register file //83-81h
		.ram_addr(a_ram_executor), //drives output RAM address (if executor control selected)
		.ram_data(d_ram_drv),		//driven by output RAM
		.selected_bit(gpi[34:32]),	//outputs address of selected bit of RAM data
		.bit_data(gpi[36]),			//outputs selected bit data
		//.tdo_1(tdo1),
		//.tdo_2(tdo2),
		//.tms_1(tms1),
		//.tms_2(tms2),
		//.tck_1(tck1),
		//.tck_2(tck2),
		.clk_cpu(clk_cpu),
		.clk_tap(clk_cpu),		//CS: drive clk_tap via on board osc and prescaler
		.mode(gpo[39:32]),	//84h
		.exec_state(gpi[47:40]),  //89h
		.run(run),
		.debug(gpi[55:48])
	);
	assign gpi[31:8] = a_ram_executor;	//for debugging executor 87-85h
	assign gpi[39:37] = 3'b000;
	assign gpi[35] = 1'b0;

	// output RAM signal mapping begin
	assign a_ram = addr_by_rf_or_ex ? gpo[31:8] : a_ram_executor; // gpo[31:8] -> 83-81h
	assign gpi[7:0] = d_ram_drv;   //read from 80h
	
		//assign d_cpu = read_en[1] ? 8'hzz : general_purpose_out [15:8];
	assign d_ram_drv = data_write_strobe ? 8'hzz : gpo[7:0];  //write to 80h	

	assign oe_ram_drv = (addr_by_rf_or_ex & data_read_strobe);
	assign wr_ram_drv_exp_mask = data_write_strobe;
	reg cs_ram;
	always @*	// make CS signal
		begin
			if (a_ram <= ram_top) cs_ram <= 1'b0;
			else cs_ram <= 1'b1;
		end
	// output RAM signal mapping end		
		
	//ram_address_manager am_out_ram (
		//.data(d_ram_drv);
	//	.addr_out(gpi[23:0]),  		// 24 bit
	//	.addr_in(gpo[31:8]),   		// 83-81h
	//	.ld_addr(addr_wrstrb),		// preload out_ram_address_manager
	//	.inc_addr(data_wrstrb),		  // L on write to 80h
	//	.reset(reset_cpu),
	//	.clk(clk_cpu),
	//	.debug(debug)
	//);
	// output RAM manager end
	



	//assign gpio_b[2] = !(command[0] | command[1]| command[2]);  // blue
	//assign gpio_b[2] = data_rd_or_wrstrb;
	//assign gpio_b[2] = data_rdstrb;
	assign gpio_b[2] = run; // blue LED on
	assign gpio_b[1] = addr_by_rf_or_ex;	// yellow LED on when exector active
	// turn blue led on in tlr or rti
	//assign gpio_b[2] = !((state == tlr) | (state == rti));
	
endmodule
